../../lab2/part1/simple_counter/simple_counter.srcs/sources_1/imports/mit6.111/binary_to_seven_seg.sv