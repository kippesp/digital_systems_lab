../../lab2/part1/simple_counter/simple_counter.srcs/sources_1/new/seven_seg_controller.sv